/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
class maxmult_sequence extends uvm_sequence #(sequence_item);
    `uvm_object_utils(maxmult_sequence)
    
//------------------------------------------------------------------------------
// local variables
//------------------------------------------------------------------------------
// not necessary, req is inherited
//    add_sequence_item req;

//------------------------------------------------------------------------------
// constructor
//------------------------------------------------------------------------------
    function new(string name = "maxmult_sequence");
        super.new(name);
    endfunction : new

//------------------------------------------------------------------------------
// the sequence body
//------------------------------------------------------------------------------
    task body();
        `uvm_info("SEQ_MIN_MAX", "", UVM_MEDIUM)
        
        `uvm_create(req);
        repeat (1000) begin
//            req = add_sequence_item::type_id::create("req");
//            start_item(req);
//            assert(req.randomize());
//            finish_item(req);
            `uvm_rand_send_with(req, {
			    arg_a dist {16'sh8000:=1, 16'sh7FFF:=1};
		        arg_b dist {16'sh8000:=1, 16'sh7FFF:=1};
			});
//            req.print();
        end
        req.rst_n = 1;
        //req.flag_arg_a_parity = 1'b0;
        //req.flag_arg_b_parity = 1'b1;
        `uvm_rand_send(req)
    endtask : body
    
    
endclass : maxmult_sequence